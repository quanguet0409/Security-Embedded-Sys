
`include "dump_file_agent.svh"
`include "csv_file_dump.svh"
`include "sample_agent.svh"
`include "loop_sample_agent.svh"
`include "sample_manager.svh"
`include "nodf_module_interface.svh"
`include "nodf_module_monitor.svh"
`include "pp_loop_interface.svh"
`include "pp_loop_monitor.svh"
`include "seq_loop_interface.svh"
`include "seq_loop_monitor.svh"
`include "upc_loop_interface.svh"
`include "upc_loop_monitor.svh"
`timescale 1ns/1ps

// top module for dataflow related monitors
module dataflow_monitor(
input logic clock,
input logic reset,
input logic finish
);



    nodf_module_intf module_intf_1(clock,reset);
    assign module_intf_1.ap_start = AESL_inst_dut.ap_start;
    assign module_intf_1.ap_ready = AESL_inst_dut.ap_ready;
    assign module_intf_1.ap_done = AESL_inst_dut.ap_done;
    assign module_intf_1.ap_continue = 1'b1;
    assign module_intf_1.finish = finish;
    csv_file_dump mstatus_csv_dumper_1;
    nodf_module_monitor module_monitor_1;
    nodf_module_intf module_intf_2(clock,reset);
    assign module_intf_2.ap_start = AESL_inst_dut.grp_dut_Pipeline_READ_LOOP_fu_5385.ap_start;
    assign module_intf_2.ap_ready = AESL_inst_dut.grp_dut_Pipeline_READ_LOOP_fu_5385.ap_ready;
    assign module_intf_2.ap_done = AESL_inst_dut.grp_dut_Pipeline_READ_LOOP_fu_5385.ap_done;
    assign module_intf_2.ap_continue = 1'b1;
    assign module_intf_2.finish = finish;
    csv_file_dump mstatus_csv_dumper_2;
    nodf_module_monitor module_monitor_2;
    nodf_module_intf module_intf_3(clock,reset);
    assign module_intf_3.ap_start = AESL_inst_dut.grp_dut_Pipeline_READ_LOOP3_fu_5392.ap_start;
    assign module_intf_3.ap_ready = AESL_inst_dut.grp_dut_Pipeline_READ_LOOP3_fu_5392.ap_ready;
    assign module_intf_3.ap_done = AESL_inst_dut.grp_dut_Pipeline_READ_LOOP3_fu_5392.ap_done;
    assign module_intf_3.ap_continue = 1'b1;
    assign module_intf_3.finish = finish;
    csv_file_dump mstatus_csv_dumper_3;
    nodf_module_monitor module_monitor_3;
    nodf_module_intf module_intf_4(clock,reset);
    assign module_intf_4.ap_start = AESL_inst_dut.grp_dut_Pipeline_READ_LOOP4_fu_5399.ap_start;
    assign module_intf_4.ap_ready = AESL_inst_dut.grp_dut_Pipeline_READ_LOOP4_fu_5399.ap_ready;
    assign module_intf_4.ap_done = AESL_inst_dut.grp_dut_Pipeline_READ_LOOP4_fu_5399.ap_done;
    assign module_intf_4.ap_continue = 1'b1;
    assign module_intf_4.finish = finish;
    csv_file_dump mstatus_csv_dumper_4;
    nodf_module_monitor module_monitor_4;
    nodf_module_intf module_intf_5(clock,reset);
    assign module_intf_5.ap_start = AESL_inst_dut.grp_dut_Pipeline_VITIS_LOOP_14_1_fu_5406.ap_start;
    assign module_intf_5.ap_ready = AESL_inst_dut.grp_dut_Pipeline_VITIS_LOOP_14_1_fu_5406.ap_ready;
    assign module_intf_5.ap_done = AESL_inst_dut.grp_dut_Pipeline_VITIS_LOOP_14_1_fu_5406.ap_done;
    assign module_intf_5.ap_continue = 1'b1;
    assign module_intf_5.finish = finish;
    csv_file_dump mstatus_csv_dumper_5;
    nodf_module_monitor module_monitor_5;
    nodf_module_intf module_intf_6(clock,reset);
    assign module_intf_6.ap_start = AESL_inst_dut.grp_divide_fu_5412.ap_start;
    assign module_intf_6.ap_ready = AESL_inst_dut.grp_divide_fu_5412.ap_ready;
    assign module_intf_6.ap_done = AESL_inst_dut.grp_divide_fu_5412.ap_done;
    assign module_intf_6.ap_continue = 1'b1;
    assign module_intf_6.finish = finish;
    csv_file_dump mstatus_csv_dumper_6;
    nodf_module_monitor module_monitor_6;
    nodf_module_intf module_intf_7(clock,reset);
    assign module_intf_7.ap_start = AESL_inst_dut.grp_divide_fu_5412.grp_divide_Pipeline_NORMALIZE_fu_2815.ap_start;
    assign module_intf_7.ap_ready = AESL_inst_dut.grp_divide_fu_5412.grp_divide_Pipeline_NORMALIZE_fu_2815.ap_ready;
    assign module_intf_7.ap_done = AESL_inst_dut.grp_divide_fu_5412.grp_divide_Pipeline_NORMALIZE_fu_2815.ap_done;
    assign module_intf_7.ap_continue = 1'b1;
    assign module_intf_7.finish = finish;
    csv_file_dump mstatus_csv_dumper_7;
    nodf_module_monitor module_monitor_7;
    nodf_module_intf module_intf_8(clock,reset);
    assign module_intf_8.ap_start = AESL_inst_dut.grp_divide_fu_5412.grp_divide_Pipeline_SHIFT_fu_2822.ap_start;
    assign module_intf_8.ap_ready = AESL_inst_dut.grp_divide_fu_5412.grp_divide_Pipeline_SHIFT_fu_2822.ap_ready;
    assign module_intf_8.ap_done = AESL_inst_dut.grp_divide_fu_5412.grp_divide_Pipeline_SHIFT_fu_2822.ap_done;
    assign module_intf_8.ap_continue = 1'b1;
    assign module_intf_8.finish = finish;
    csv_file_dump mstatus_csv_dumper_8;
    nodf_module_monitor module_monitor_8;
    nodf_module_intf module_intf_9(clock,reset);
    assign module_intf_9.ap_start = AESL_inst_dut.grp_divide_fu_5412.grp_divide_Pipeline_SHIFT5_fu_2838.ap_start;
    assign module_intf_9.ap_ready = AESL_inst_dut.grp_divide_fu_5412.grp_divide_Pipeline_SHIFT5_fu_2838.ap_ready;
    assign module_intf_9.ap_done = AESL_inst_dut.grp_divide_fu_5412.grp_divide_Pipeline_SHIFT5_fu_2838.ap_done;
    assign module_intf_9.ap_continue = 1'b1;
    assign module_intf_9.finish = finish;
    csv_file_dump mstatus_csv_dumper_9;
    nodf_module_monitor module_monitor_9;
    nodf_module_intf module_intf_10(clock,reset);
    assign module_intf_10.ap_start = AESL_inst_dut.grp_divide_fu_5412.grp_divide_Pipeline_CLEAR_UPPER_fu_2854.ap_start;
    assign module_intf_10.ap_ready = AESL_inst_dut.grp_divide_fu_5412.grp_divide_Pipeline_CLEAR_UPPER_fu_2854.ap_ready;
    assign module_intf_10.ap_done = AESL_inst_dut.grp_divide_fu_5412.grp_divide_Pipeline_CLEAR_UPPER_fu_2854.ap_done;
    assign module_intf_10.ap_continue = 1'b1;
    assign module_intf_10.finish = finish;
    csv_file_dump mstatus_csv_dumper_10;
    nodf_module_monitor module_monitor_10;
    nodf_module_intf module_intf_11(clock,reset);
    assign module_intf_11.ap_start = AESL_inst_dut.grp_divide_fu_5412.grp_divide_Pipeline_PARTIAL_fu_2864.ap_start;
    assign module_intf_11.ap_ready = AESL_inst_dut.grp_divide_fu_5412.grp_divide_Pipeline_PARTIAL_fu_2864.ap_ready;
    assign module_intf_11.ap_done = AESL_inst_dut.grp_divide_fu_5412.grp_divide_Pipeline_PARTIAL_fu_2864.ap_done;
    assign module_intf_11.ap_continue = 1'b1;
    assign module_intf_11.finish = finish;
    csv_file_dump mstatus_csv_dumper_11;
    nodf_module_monitor module_monitor_11;
    nodf_module_intf module_intf_12(clock,reset);
    assign module_intf_12.ap_start = AESL_inst_dut.grp_divide_fu_5412.grp_divide_Pipeline_COMPARE_fu_2878.ap_start;
    assign module_intf_12.ap_ready = AESL_inst_dut.grp_divide_fu_5412.grp_divide_Pipeline_COMPARE_fu_2878.ap_ready;
    assign module_intf_12.ap_done = AESL_inst_dut.grp_divide_fu_5412.grp_divide_Pipeline_COMPARE_fu_2878.ap_done;
    assign module_intf_12.ap_continue = 1'b1;
    assign module_intf_12.finish = finish;
    csv_file_dump mstatus_csv_dumper_12;
    nodf_module_monitor module_monitor_12;
    nodf_module_intf module_intf_13(clock,reset);
    assign module_intf_13.ap_start = AESL_inst_dut.grp_divide_fu_5412.grp_divide_Pipeline_ADJUST_fu_2889.ap_start;
    assign module_intf_13.ap_ready = AESL_inst_dut.grp_divide_fu_5412.grp_divide_Pipeline_ADJUST_fu_2889.ap_ready;
    assign module_intf_13.ap_done = AESL_inst_dut.grp_divide_fu_5412.grp_divide_Pipeline_ADJUST_fu_2889.ap_done;
    assign module_intf_13.ap_continue = 1'b1;
    assign module_intf_13.finish = finish;
    csv_file_dump mstatus_csv_dumper_13;
    nodf_module_monitor module_monitor_13;
    nodf_module_intf module_intf_14(clock,reset);
    assign module_intf_14.ap_start = AESL_inst_dut.grp_divide_fu_5412.grp_divide_Pipeline_REM_fu_2899.ap_start;
    assign module_intf_14.ap_ready = AESL_inst_dut.grp_divide_fu_5412.grp_divide_Pipeline_REM_fu_2899.ap_ready;
    assign module_intf_14.ap_done = AESL_inst_dut.grp_divide_fu_5412.grp_divide_Pipeline_REM_fu_2899.ap_done;
    assign module_intf_14.ap_continue = 1'b1;
    assign module_intf_14.finish = finish;
    csv_file_dump mstatus_csv_dumper_14;
    nodf_module_monitor module_monitor_14;
    nodf_module_intf module_intf_15(clock,reset);
    assign module_intf_15.ap_start = AESL_inst_dut.grp_divide_fu_5412.grp_divide_Pipeline_SHIFT6_fu_2911.ap_start;
    assign module_intf_15.ap_ready = AESL_inst_dut.grp_divide_fu_5412.grp_divide_Pipeline_SHIFT6_fu_2911.ap_ready;
    assign module_intf_15.ap_done = AESL_inst_dut.grp_divide_fu_5412.grp_divide_Pipeline_SHIFT6_fu_2911.ap_done;
    assign module_intf_15.ap_continue = 1'b1;
    assign module_intf_15.finish = finish;
    csv_file_dump mstatus_csv_dumper_15;
    nodf_module_monitor module_monitor_15;
    nodf_module_intf module_intf_16(clock,reset);
    assign module_intf_16.ap_start = AESL_inst_dut.grp_operator_lt_fu_5420.ap_start;
    assign module_intf_16.ap_ready = AESL_inst_dut.grp_operator_lt_fu_5420.ap_ready;
    assign module_intf_16.ap_done = AESL_inst_dut.grp_operator_lt_fu_5420.ap_done;
    assign module_intf_16.ap_continue = 1'b1;
    assign module_intf_16.finish = finish;
    csv_file_dump mstatus_csv_dumper_16;
    nodf_module_monitor module_monitor_16;
    nodf_module_intf module_intf_17(clock,reset);
    assign module_intf_17.ap_start = AESL_inst_dut.grp_operator_mul_fu_5426.ap_start;
    assign module_intf_17.ap_ready = AESL_inst_dut.grp_operator_mul_fu_5426.ap_ready;
    assign module_intf_17.ap_done = AESL_inst_dut.grp_operator_mul_fu_5426.ap_done;
    assign module_intf_17.ap_continue = 1'b1;
    assign module_intf_17.finish = finish;
    csv_file_dump mstatus_csv_dumper_17;
    nodf_module_monitor module_monitor_17;
    nodf_module_intf module_intf_18(clock,reset);
    assign module_intf_18.ap_start = AESL_inst_dut.grp_operator_mul_fu_5426.grp_operator_Pipeline_OUTER_INNER_fu_371.ap_start;
    assign module_intf_18.ap_ready = AESL_inst_dut.grp_operator_mul_fu_5426.grp_operator_Pipeline_OUTER_INNER_fu_371.ap_ready;
    assign module_intf_18.ap_done = AESL_inst_dut.grp_operator_mul_fu_5426.grp_operator_Pipeline_OUTER_INNER_fu_371.ap_done;
    assign module_intf_18.ap_continue = 1'b1;
    assign module_intf_18.finish = finish;
    csv_file_dump mstatus_csv_dumper_18;
    nodf_module_monitor module_monitor_18;
    nodf_module_intf module_intf_19(clock,reset);
    assign module_intf_19.ap_start = AESL_inst_dut.grp_dut_Pipeline_SHIFT_fu_5433.ap_start;
    assign module_intf_19.ap_ready = AESL_inst_dut.grp_dut_Pipeline_SHIFT_fu_5433.ap_ready;
    assign module_intf_19.ap_done = AESL_inst_dut.grp_dut_Pipeline_SHIFT_fu_5433.ap_done;
    assign module_intf_19.ap_continue = 1'b1;
    assign module_intf_19.finish = finish;
    csv_file_dump mstatus_csv_dumper_19;
    nodf_module_monitor module_monitor_19;
    nodf_module_intf module_intf_20(clock,reset);
    assign module_intf_20.ap_start = AESL_inst_dut.grp_operator_1_fu_5440.ap_start;
    assign module_intf_20.ap_ready = AESL_inst_dut.grp_operator_1_fu_5440.ap_ready;
    assign module_intf_20.ap_done = AESL_inst_dut.grp_operator_1_fu_5440.ap_done;
    assign module_intf_20.ap_continue = 1'b1;
    assign module_intf_20.finish = finish;
    csv_file_dump mstatus_csv_dumper_20;
    nodf_module_monitor module_monitor_20;
    nodf_module_intf module_intf_21(clock,reset);
    assign module_intf_21.ap_start = AESL_inst_dut.grp_operator_1_fu_5440.grp_operator_1_Pipeline_OUTER_INNER_fu_369.ap_start;
    assign module_intf_21.ap_ready = AESL_inst_dut.grp_operator_1_fu_5440.grp_operator_1_Pipeline_OUTER_INNER_fu_369.ap_ready;
    assign module_intf_21.ap_done = AESL_inst_dut.grp_operator_1_fu_5440.grp_operator_1_Pipeline_OUTER_INNER_fu_369.ap_done;
    assign module_intf_21.ap_continue = 1'b1;
    assign module_intf_21.finish = finish;
    csv_file_dump mstatus_csv_dumper_21;
    nodf_module_monitor module_monitor_21;
    nodf_module_intf module_intf_22(clock,reset);
    assign module_intf_22.ap_start = AESL_inst_dut.grp_dut_Pipeline_WRITE_LOOP_fu_5446.ap_start;
    assign module_intf_22.ap_ready = AESL_inst_dut.grp_dut_Pipeline_WRITE_LOOP_fu_5446.ap_ready;
    assign module_intf_22.ap_done = AESL_inst_dut.grp_dut_Pipeline_WRITE_LOOP_fu_5446.ap_done;
    assign module_intf_22.ap_continue = 1'b1;
    assign module_intf_22.finish = finish;
    csv_file_dump mstatus_csv_dumper_22;
    nodf_module_monitor module_monitor_22;

    pp_loop_intf #(7) pp_loop_intf_1(clock,reset);
    assign pp_loop_intf_1.pre_loop_state0 = AESL_inst_dut.grp_divide_fu_5412.grp_divide_Pipeline_SHIFT_fu_2822.ap_ST_fsm_state1;
    assign pp_loop_intf_1.pre_states_valid = 1'b1;
    assign pp_loop_intf_1.post_loop_state0 = AESL_inst_dut.grp_divide_fu_5412.grp_divide_Pipeline_SHIFT_fu_2822.ap_ST_fsm_state8;
    assign pp_loop_intf_1.post_states_valid[0] = 1'b1;
    assign pp_loop_intf_1.post_loop_state1 = AESL_inst_dut.grp_divide_fu_5412.grp_divide_Pipeline_SHIFT_fu_2822.ap_ST_fsm_state9;
    assign pp_loop_intf_1.post_states_valid[1] = 1'b1;
    assign pp_loop_intf_1.post_loop_state2 = AESL_inst_dut.grp_divide_fu_5412.grp_divide_Pipeline_SHIFT_fu_2822.ap_ST_fsm_state10;
    assign pp_loop_intf_1.post_states_valid[2] = 1'b1;
    assign pp_loop_intf_1.iter_start_state = AESL_inst_dut.grp_divide_fu_5412.grp_divide_Pipeline_SHIFT_fu_2822.ap_ST_fsm_pp0_stage0;
    assign pp_loop_intf_1.iter_start_enable = AESL_inst_dut.grp_divide_fu_5412.grp_divide_Pipeline_SHIFT_fu_2822.ap_enable_reg_pp0_iter0;
    assign pp_loop_intf_1.iter_start_block = AESL_inst_dut.grp_divide_fu_5412.grp_divide_Pipeline_SHIFT_fu_2822.ap_block_pp0_stage0_subdone;
    assign pp_loop_intf_1.iter_end_state = AESL_inst_dut.grp_divide_fu_5412.grp_divide_Pipeline_SHIFT_fu_2822.ap_ST_fsm_pp0_stage1;
    assign pp_loop_intf_1.iter_end_enable = AESL_inst_dut.grp_divide_fu_5412.grp_divide_Pipeline_SHIFT_fu_2822.ap_enable_reg_pp0_iter2;
    assign pp_loop_intf_1.iter_end_block = AESL_inst_dut.grp_divide_fu_5412.grp_divide_Pipeline_SHIFT_fu_2822.ap_block_pp0_stage1_subdone;
    assign pp_loop_intf_1.loop_quit_state = AESL_inst_dut.grp_divide_fu_5412.grp_divide_Pipeline_SHIFT_fu_2822.ap_ST_fsm_pp0_stage1;
    assign pp_loop_intf_1.quit_at_end = 1'b0;
    assign pp_loop_intf_1.cur_state = AESL_inst_dut.grp_divide_fu_5412.grp_divide_Pipeline_SHIFT_fu_2822.ap_CS_fsm;
    assign pp_loop_intf_1.finish = finish;
    csv_file_dump pp_loop_csv_dumper_1;
    pp_loop_monitor #(7) pp_loop_monitor_1;
    pp_loop_intf #(7) pp_loop_intf_2(clock,reset);
    assign pp_loop_intf_2.pre_loop_state0 = AESL_inst_dut.grp_divide_fu_5412.grp_divide_Pipeline_SHIFT5_fu_2838.ap_ST_fsm_state1;
    assign pp_loop_intf_2.pre_states_valid = 1'b1;
    assign pp_loop_intf_2.post_loop_state0 = AESL_inst_dut.grp_divide_fu_5412.grp_divide_Pipeline_SHIFT5_fu_2838.ap_ST_fsm_state8;
    assign pp_loop_intf_2.post_states_valid[0] = 1'b1;
    assign pp_loop_intf_2.post_loop_state1 = AESL_inst_dut.grp_divide_fu_5412.grp_divide_Pipeline_SHIFT5_fu_2838.ap_ST_fsm_state9;
    assign pp_loop_intf_2.post_states_valid[1] = 1'b1;
    assign pp_loop_intf_2.post_loop_state2 = AESL_inst_dut.grp_divide_fu_5412.grp_divide_Pipeline_SHIFT5_fu_2838.ap_ST_fsm_state10;
    assign pp_loop_intf_2.post_states_valid[2] = 1'b1;
    assign pp_loop_intf_2.iter_start_state = AESL_inst_dut.grp_divide_fu_5412.grp_divide_Pipeline_SHIFT5_fu_2838.ap_ST_fsm_pp0_stage0;
    assign pp_loop_intf_2.iter_start_enable = AESL_inst_dut.grp_divide_fu_5412.grp_divide_Pipeline_SHIFT5_fu_2838.ap_enable_reg_pp0_iter0;
    assign pp_loop_intf_2.iter_start_block = AESL_inst_dut.grp_divide_fu_5412.grp_divide_Pipeline_SHIFT5_fu_2838.ap_block_pp0_stage0_subdone;
    assign pp_loop_intf_2.iter_end_state = AESL_inst_dut.grp_divide_fu_5412.grp_divide_Pipeline_SHIFT5_fu_2838.ap_ST_fsm_pp0_stage1;
    assign pp_loop_intf_2.iter_end_enable = AESL_inst_dut.grp_divide_fu_5412.grp_divide_Pipeline_SHIFT5_fu_2838.ap_enable_reg_pp0_iter2;
    assign pp_loop_intf_2.iter_end_block = AESL_inst_dut.grp_divide_fu_5412.grp_divide_Pipeline_SHIFT5_fu_2838.ap_block_pp0_stage1_subdone;
    assign pp_loop_intf_2.loop_quit_state = AESL_inst_dut.grp_divide_fu_5412.grp_divide_Pipeline_SHIFT5_fu_2838.ap_ST_fsm_pp0_stage1;
    assign pp_loop_intf_2.quit_at_end = 1'b0;
    assign pp_loop_intf_2.cur_state = AESL_inst_dut.grp_divide_fu_5412.grp_divide_Pipeline_SHIFT5_fu_2838.ap_CS_fsm;
    assign pp_loop_intf_2.finish = finish;
    csv_file_dump pp_loop_csv_dumper_2;
    pp_loop_monitor #(7) pp_loop_monitor_2;
    pp_loop_intf #(6) pp_loop_intf_3(clock,reset);
    assign pp_loop_intf_3.pre_loop_state0 = AESL_inst_dut.grp_divide_fu_5412.grp_divide_Pipeline_PARTIAL_fu_2864.ap_ST_fsm_state1;
    assign pp_loop_intf_3.pre_states_valid = 1'b1;
    assign pp_loop_intf_3.post_loop_state0 = AESL_inst_dut.grp_divide_fu_5412.grp_divide_Pipeline_PARTIAL_fu_2864.ap_ST_fsm_state10;
    assign pp_loop_intf_3.post_states_valid[0] = 1'b1;
    assign pp_loop_intf_3.post_loop_state1 = AESL_inst_dut.grp_divide_fu_5412.grp_divide_Pipeline_PARTIAL_fu_2864.ap_ST_fsm_state11;
    assign pp_loop_intf_3.post_states_valid[1] = 1'b1;
    assign pp_loop_intf_3.post_loop_state2 = AESL_inst_dut.grp_divide_fu_5412.grp_divide_Pipeline_PARTIAL_fu_2864.ap_ST_fsm_state12;
    assign pp_loop_intf_3.post_states_valid[2] = 1'b1;
    assign pp_loop_intf_3.iter_start_state = AESL_inst_dut.grp_divide_fu_5412.grp_divide_Pipeline_PARTIAL_fu_2864.ap_ST_fsm_pp0_stage0;
    assign pp_loop_intf_3.iter_start_enable = AESL_inst_dut.grp_divide_fu_5412.grp_divide_Pipeline_PARTIAL_fu_2864.ap_enable_reg_pp0_iter0;
    assign pp_loop_intf_3.iter_start_block = AESL_inst_dut.grp_divide_fu_5412.grp_divide_Pipeline_PARTIAL_fu_2864.ap_block_pp0_stage0_subdone;
    assign pp_loop_intf_3.iter_end_state = AESL_inst_dut.grp_divide_fu_5412.grp_divide_Pipeline_PARTIAL_fu_2864.ap_ST_fsm_pp0_stage1;
    assign pp_loop_intf_3.iter_end_enable = AESL_inst_dut.grp_divide_fu_5412.grp_divide_Pipeline_PARTIAL_fu_2864.ap_enable_reg_pp0_iter3;
    assign pp_loop_intf_3.iter_end_block = AESL_inst_dut.grp_divide_fu_5412.grp_divide_Pipeline_PARTIAL_fu_2864.ap_block_pp0_stage1_subdone;
    assign pp_loop_intf_3.loop_quit_state = AESL_inst_dut.grp_divide_fu_5412.grp_divide_Pipeline_PARTIAL_fu_2864.ap_ST_fsm_pp0_stage0;
    assign pp_loop_intf_3.quit_at_end = 1'b0;
    assign pp_loop_intf_3.cur_state = AESL_inst_dut.grp_divide_fu_5412.grp_divide_Pipeline_PARTIAL_fu_2864.ap_CS_fsm;
    assign pp_loop_intf_3.finish = finish;
    csv_file_dump pp_loop_csv_dumper_3;
    pp_loop_monitor #(6) pp_loop_monitor_3;
    seq_loop_intf#(251) seq_loop_intf_1(clock,reset);
    assign seq_loop_intf_1.pre_loop_state0 = AESL_inst_dut.ap_ST_fsm_state79;
    assign seq_loop_intf_1.pre_states_valid = 1'b1;
    assign seq_loop_intf_1.post_loop_state0 = AESL_inst_dut.ap_ST_fsm_state218;
    assign seq_loop_intf_1.post_states_valid[0] = 1'b1;
    assign seq_loop_intf_1.post_loop_state1 = 251'h0;
    assign seq_loop_intf_1.post_states_valid[1] = 1'b0;
    assign seq_loop_intf_1.post_loop_state2 = 251'h0;
    assign seq_loop_intf_1.post_states_valid[2] = 1'b0;
    assign seq_loop_intf_1.post_loop_state3 = 251'h0;
    assign seq_loop_intf_1.post_states_valid[3] = 1'b0;
    assign seq_loop_intf_1.post_loop_state4 = 251'h0;
    assign seq_loop_intf_1.post_states_valid[4] = 1'b0;
    assign seq_loop_intf_1.quit_loop_state0 = AESL_inst_dut.ap_ST_fsm_state80;
    assign seq_loop_intf_1.quit_states_valid = 1'b1;
    assign seq_loop_intf_1.cur_state = AESL_inst_dut.ap_CS_fsm;
    assign seq_loop_intf_1.iter_start_state = AESL_inst_dut.ap_ST_fsm_state80;
    assign seq_loop_intf_1.iter_end_state0 = AESL_inst_dut.ap_ST_fsm_state217;
    assign seq_loop_intf_1.iter_end_states_valid = 1'b1;
    assign seq_loop_intf_1.one_state_loop = 1'b0;
    assign seq_loop_intf_1.one_state_block = 1'b0;
    assign seq_loop_intf_1.finish = finish;
    csv_file_dump seq_loop_csv_dumper_1;
    seq_loop_monitor #(251) seq_loop_monitor_1;
    seq_loop_intf#(459) seq_loop_intf_2(clock,reset);
    assign seq_loop_intf_2.pre_loop_state0 = AESL_inst_dut.grp_divide_fu_5412.ap_ST_fsm_state81;
    assign seq_loop_intf_2.pre_states_valid = 1'b1;
    assign seq_loop_intf_2.post_loop_state0 = AESL_inst_dut.grp_divide_fu_5412.ap_ST_fsm_state84;
    assign seq_loop_intf_2.post_states_valid[0] = 1'b1;
    assign seq_loop_intf_2.post_loop_state1 = AESL_inst_dut.grp_divide_fu_5412.ap_ST_fsm_state83;
    assign seq_loop_intf_2.post_states_valid[1] = 1'b1;
    assign seq_loop_intf_2.post_loop_state2 = 459'h0;
    assign seq_loop_intf_2.post_states_valid[2] = 1'b0;
    assign seq_loop_intf_2.post_loop_state3 = 459'h0;
    assign seq_loop_intf_2.post_states_valid[3] = 1'b0;
    assign seq_loop_intf_2.post_loop_state4 = 459'h0;
    assign seq_loop_intf_2.post_states_valid[4] = 1'b0;
    assign seq_loop_intf_2.quit_loop_state0 = AESL_inst_dut.grp_divide_fu_5412.ap_ST_fsm_state82;
    assign seq_loop_intf_2.quit_states_valid = 1'b1;
    assign seq_loop_intf_2.cur_state = AESL_inst_dut.grp_divide_fu_5412.ap_CS_fsm;
    assign seq_loop_intf_2.iter_start_state = AESL_inst_dut.grp_divide_fu_5412.ap_ST_fsm_state82;
    assign seq_loop_intf_2.iter_end_state0 = AESL_inst_dut.grp_divide_fu_5412.ap_ST_fsm_state82;
    assign seq_loop_intf_2.iter_end_states_valid = 1'b1;
    assign seq_loop_intf_2.one_state_loop = 1'b1;
    assign seq_loop_intf_2.one_state_block = AESL_inst_dut.grp_divide_fu_5412.ap_ST_fsm_state82_blk;
    assign seq_loop_intf_2.finish = finish;
    csv_file_dump seq_loop_csv_dumper_2;
    seq_loop_monitor #(459) seq_loop_monitor_2;
    seq_loop_intf#(459) seq_loop_intf_3(clock,reset);
    assign seq_loop_intf_3.pre_loop_state0 = AESL_inst_dut.grp_divide_fu_5412.ap_ST_fsm_state381;
    assign seq_loop_intf_3.pre_states_valid = 1'b1;
    assign seq_loop_intf_3.post_loop_state0 = AESL_inst_dut.grp_divide_fu_5412.ap_ST_fsm_state393;
    assign seq_loop_intf_3.post_states_valid[0] = 1'b1;
    assign seq_loop_intf_3.post_loop_state1 = 459'h0;
    assign seq_loop_intf_3.post_states_valid[1] = 1'b0;
    assign seq_loop_intf_3.post_loop_state2 = 459'h0;
    assign seq_loop_intf_3.post_states_valid[2] = 1'b0;
    assign seq_loop_intf_3.post_loop_state3 = 459'h0;
    assign seq_loop_intf_3.post_states_valid[3] = 1'b0;
    assign seq_loop_intf_3.post_loop_state4 = 459'h0;
    assign seq_loop_intf_3.post_states_valid[4] = 1'b0;
    assign seq_loop_intf_3.quit_loop_state0 = AESL_inst_dut.grp_divide_fu_5412.ap_ST_fsm_state386;
    assign seq_loop_intf_3.quit_states_valid = 1'b1;
    assign seq_loop_intf_3.cur_state = AESL_inst_dut.grp_divide_fu_5412.ap_CS_fsm;
    assign seq_loop_intf_3.iter_start_state = AESL_inst_dut.grp_divide_fu_5412.ap_ST_fsm_state382;
    assign seq_loop_intf_3.iter_end_state0 = AESL_inst_dut.grp_divide_fu_5412.ap_ST_fsm_state392;
    assign seq_loop_intf_3.iter_end_states_valid = 1'b1;
    assign seq_loop_intf_3.one_state_loop = 1'b0;
    assign seq_loop_intf_3.one_state_block = 1'b0;
    assign seq_loop_intf_3.finish = finish;
    csv_file_dump seq_loop_csv_dumper_3;
    seq_loop_monitor #(459) seq_loop_monitor_3;
    seq_loop_intf#(459) seq_loop_intf_4(clock,reset);
    assign seq_loop_intf_4.pre_loop_state0 = AESL_inst_dut.grp_divide_fu_5412.ap_ST_fsm_state243;
    assign seq_loop_intf_4.pre_states_valid = 1'b1;
    assign seq_loop_intf_4.post_loop_state0 = AESL_inst_dut.grp_divide_fu_5412.ap_ST_fsm_state395;
    assign seq_loop_intf_4.post_states_valid[0] = 1'b1;
    assign seq_loop_intf_4.post_loop_state1 = 459'h0;
    assign seq_loop_intf_4.post_states_valid[1] = 1'b0;
    assign seq_loop_intf_4.post_loop_state2 = 459'h0;
    assign seq_loop_intf_4.post_states_valid[2] = 1'b0;
    assign seq_loop_intf_4.post_loop_state3 = 459'h0;
    assign seq_loop_intf_4.post_states_valid[3] = 1'b0;
    assign seq_loop_intf_4.post_loop_state4 = 459'h0;
    assign seq_loop_intf_4.post_states_valid[4] = 1'b0;
    assign seq_loop_intf_4.quit_loop_state0 = AESL_inst_dut.grp_divide_fu_5412.ap_ST_fsm_state244;
    assign seq_loop_intf_4.quit_states_valid = 1'b1;
    assign seq_loop_intf_4.cur_state = AESL_inst_dut.grp_divide_fu_5412.ap_CS_fsm;
    assign seq_loop_intf_4.iter_start_state = AESL_inst_dut.grp_divide_fu_5412.ap_ST_fsm_state244;
    assign seq_loop_intf_4.iter_end_state0 = AESL_inst_dut.grp_divide_fu_5412.ap_ST_fsm_state394;
    assign seq_loop_intf_4.iter_end_states_valid = 1'b1;
    assign seq_loop_intf_4.one_state_loop = 1'b0;
    assign seq_loop_intf_4.one_state_block = 1'b0;
    assign seq_loop_intf_4.finish = finish;
    csv_file_dump seq_loop_csv_dumper_4;
    seq_loop_monitor #(459) seq_loop_monitor_4;
    seq_loop_intf#(12) seq_loop_intf_5(clock,reset);
    assign seq_loop_intf_5.pre_loop_state0 = AESL_inst_dut.grp_divide_fu_5412.grp_divide_Pipeline_COMPARE_fu_2878.ap_ST_fsm_state1;
    assign seq_loop_intf_5.pre_states_valid = 1'b1;
    assign seq_loop_intf_5.post_loop_state0 = AESL_inst_dut.grp_divide_fu_5412.grp_divide_Pipeline_COMPARE_fu_2878.ap_ST_fsm_state8;
    assign seq_loop_intf_5.post_states_valid[0] = 1'b1;
    assign seq_loop_intf_5.post_loop_state1 = AESL_inst_dut.grp_divide_fu_5412.grp_divide_Pipeline_COMPARE_fu_2878.ap_ST_fsm_state9;
    assign seq_loop_intf_5.post_states_valid[1] = 1'b1;
    assign seq_loop_intf_5.post_loop_state2 = AESL_inst_dut.grp_divide_fu_5412.grp_divide_Pipeline_COMPARE_fu_2878.ap_ST_fsm_state10;
    assign seq_loop_intf_5.post_states_valid[2] = 1'b1;
    assign seq_loop_intf_5.post_loop_state3 = AESL_inst_dut.grp_divide_fu_5412.grp_divide_Pipeline_COMPARE_fu_2878.ap_ST_fsm_state11;
    assign seq_loop_intf_5.post_states_valid[3] = 1'b1;
    assign seq_loop_intf_5.post_loop_state4 = AESL_inst_dut.grp_divide_fu_5412.grp_divide_Pipeline_COMPARE_fu_2878.ap_ST_fsm_state12;
    assign seq_loop_intf_5.post_states_valid[4] = 1'b1;
    assign seq_loop_intf_5.quit_loop_state0 = AESL_inst_dut.grp_divide_fu_5412.grp_divide_Pipeline_COMPARE_fu_2878.ap_ST_fsm_state7;
    assign seq_loop_intf_5.quit_states_valid = 1'b1;
    assign seq_loop_intf_5.cur_state = AESL_inst_dut.grp_divide_fu_5412.grp_divide_Pipeline_COMPARE_fu_2878.ap_CS_fsm;
    assign seq_loop_intf_5.iter_start_state = AESL_inst_dut.grp_divide_fu_5412.grp_divide_Pipeline_COMPARE_fu_2878.ap_ST_fsm_state2;
    assign seq_loop_intf_5.iter_end_state0 = AESL_inst_dut.grp_divide_fu_5412.grp_divide_Pipeline_COMPARE_fu_2878.ap_ST_fsm_state7;
    assign seq_loop_intf_5.iter_end_states_valid = 1'b1;
    assign seq_loop_intf_5.one_state_loop = 1'b0;
    assign seq_loop_intf_5.one_state_block = 1'b0;
    assign seq_loop_intf_5.finish = finish;
    csv_file_dump seq_loop_csv_dumper_5;
    seq_loop_monitor #(12) seq_loop_monitor_5;
    upc_loop_intf#(2) upc_loop_intf_1(clock,reset);
    assign upc_loop_intf_1.cur_state = AESL_inst_dut.grp_dut_Pipeline_READ_LOOP_fu_5385.ap_CS_fsm;
    assign upc_loop_intf_1.iter_start_state = AESL_inst_dut.grp_dut_Pipeline_READ_LOOP_fu_5385.ap_ST_fsm_pp0_stage0;
    assign upc_loop_intf_1.iter_end_state = AESL_inst_dut.grp_dut_Pipeline_READ_LOOP_fu_5385.ap_ST_fsm_pp0_stage1;
    assign upc_loop_intf_1.quit_state = AESL_inst_dut.grp_dut_Pipeline_READ_LOOP_fu_5385.ap_ST_fsm_pp0_stage1;
    assign upc_loop_intf_1.iter_start_block = AESL_inst_dut.grp_dut_Pipeline_READ_LOOP_fu_5385.ap_block_pp0_stage0_subdone;
    assign upc_loop_intf_1.iter_end_block = AESL_inst_dut.grp_dut_Pipeline_READ_LOOP_fu_5385.ap_block_pp0_stage1_subdone;
    assign upc_loop_intf_1.quit_block = AESL_inst_dut.grp_dut_Pipeline_READ_LOOP_fu_5385.ap_block_pp0_stage1_subdone;
    assign upc_loop_intf_1.iter_start_enable = AESL_inst_dut.grp_dut_Pipeline_READ_LOOP_fu_5385.ap_enable_reg_pp0_iter0;
    assign upc_loop_intf_1.iter_end_enable = AESL_inst_dut.grp_dut_Pipeline_READ_LOOP_fu_5385.ap_enable_reg_pp0_iter1;
    assign upc_loop_intf_1.quit_enable = AESL_inst_dut.grp_dut_Pipeline_READ_LOOP_fu_5385.ap_enable_reg_pp0_iter1;
    assign upc_loop_intf_1.loop_start = AESL_inst_dut.grp_dut_Pipeline_READ_LOOP_fu_5385.ap_start;
    assign upc_loop_intf_1.loop_ready = AESL_inst_dut.grp_dut_Pipeline_READ_LOOP_fu_5385.ap_ready;
    assign upc_loop_intf_1.loop_done = AESL_inst_dut.grp_dut_Pipeline_READ_LOOP_fu_5385.ap_done_int;
    assign upc_loop_intf_1.loop_continue = 1'b1;
    assign upc_loop_intf_1.quit_at_end = 1'b1;
    assign upc_loop_intf_1.finish = finish;
    csv_file_dump upc_loop_csv_dumper_1;
    upc_loop_monitor #(2) upc_loop_monitor_1;
    upc_loop_intf#(2) upc_loop_intf_2(clock,reset);
    assign upc_loop_intf_2.cur_state = AESL_inst_dut.grp_dut_Pipeline_READ_LOOP3_fu_5392.ap_CS_fsm;
    assign upc_loop_intf_2.iter_start_state = AESL_inst_dut.grp_dut_Pipeline_READ_LOOP3_fu_5392.ap_ST_fsm_pp0_stage0;
    assign upc_loop_intf_2.iter_end_state = AESL_inst_dut.grp_dut_Pipeline_READ_LOOP3_fu_5392.ap_ST_fsm_pp0_stage1;
    assign upc_loop_intf_2.quit_state = AESL_inst_dut.grp_dut_Pipeline_READ_LOOP3_fu_5392.ap_ST_fsm_pp0_stage1;
    assign upc_loop_intf_2.iter_start_block = AESL_inst_dut.grp_dut_Pipeline_READ_LOOP3_fu_5392.ap_block_pp0_stage0_subdone;
    assign upc_loop_intf_2.iter_end_block = AESL_inst_dut.grp_dut_Pipeline_READ_LOOP3_fu_5392.ap_block_pp0_stage1_subdone;
    assign upc_loop_intf_2.quit_block = AESL_inst_dut.grp_dut_Pipeline_READ_LOOP3_fu_5392.ap_block_pp0_stage1_subdone;
    assign upc_loop_intf_2.iter_start_enable = AESL_inst_dut.grp_dut_Pipeline_READ_LOOP3_fu_5392.ap_enable_reg_pp0_iter0;
    assign upc_loop_intf_2.iter_end_enable = AESL_inst_dut.grp_dut_Pipeline_READ_LOOP3_fu_5392.ap_enable_reg_pp0_iter1;
    assign upc_loop_intf_2.quit_enable = AESL_inst_dut.grp_dut_Pipeline_READ_LOOP3_fu_5392.ap_enable_reg_pp0_iter1;
    assign upc_loop_intf_2.loop_start = AESL_inst_dut.grp_dut_Pipeline_READ_LOOP3_fu_5392.ap_start;
    assign upc_loop_intf_2.loop_ready = AESL_inst_dut.grp_dut_Pipeline_READ_LOOP3_fu_5392.ap_ready;
    assign upc_loop_intf_2.loop_done = AESL_inst_dut.grp_dut_Pipeline_READ_LOOP3_fu_5392.ap_done_int;
    assign upc_loop_intf_2.loop_continue = 1'b1;
    assign upc_loop_intf_2.quit_at_end = 1'b1;
    assign upc_loop_intf_2.finish = finish;
    csv_file_dump upc_loop_csv_dumper_2;
    upc_loop_monitor #(2) upc_loop_monitor_2;
    upc_loop_intf#(2) upc_loop_intf_3(clock,reset);
    assign upc_loop_intf_3.cur_state = AESL_inst_dut.grp_dut_Pipeline_READ_LOOP4_fu_5399.ap_CS_fsm;
    assign upc_loop_intf_3.iter_start_state = AESL_inst_dut.grp_dut_Pipeline_READ_LOOP4_fu_5399.ap_ST_fsm_pp0_stage0;
    assign upc_loop_intf_3.iter_end_state = AESL_inst_dut.grp_dut_Pipeline_READ_LOOP4_fu_5399.ap_ST_fsm_pp0_stage1;
    assign upc_loop_intf_3.quit_state = AESL_inst_dut.grp_dut_Pipeline_READ_LOOP4_fu_5399.ap_ST_fsm_pp0_stage1;
    assign upc_loop_intf_3.iter_start_block = AESL_inst_dut.grp_dut_Pipeline_READ_LOOP4_fu_5399.ap_block_pp0_stage0_subdone;
    assign upc_loop_intf_3.iter_end_block = AESL_inst_dut.grp_dut_Pipeline_READ_LOOP4_fu_5399.ap_block_pp0_stage1_subdone;
    assign upc_loop_intf_3.quit_block = AESL_inst_dut.grp_dut_Pipeline_READ_LOOP4_fu_5399.ap_block_pp0_stage1_subdone;
    assign upc_loop_intf_3.iter_start_enable = AESL_inst_dut.grp_dut_Pipeline_READ_LOOP4_fu_5399.ap_enable_reg_pp0_iter0;
    assign upc_loop_intf_3.iter_end_enable = AESL_inst_dut.grp_dut_Pipeline_READ_LOOP4_fu_5399.ap_enable_reg_pp0_iter1;
    assign upc_loop_intf_3.quit_enable = AESL_inst_dut.grp_dut_Pipeline_READ_LOOP4_fu_5399.ap_enable_reg_pp0_iter1;
    assign upc_loop_intf_3.loop_start = AESL_inst_dut.grp_dut_Pipeline_READ_LOOP4_fu_5399.ap_start;
    assign upc_loop_intf_3.loop_ready = AESL_inst_dut.grp_dut_Pipeline_READ_LOOP4_fu_5399.ap_ready;
    assign upc_loop_intf_3.loop_done = AESL_inst_dut.grp_dut_Pipeline_READ_LOOP4_fu_5399.ap_done_int;
    assign upc_loop_intf_3.loop_continue = 1'b1;
    assign upc_loop_intf_3.quit_at_end = 1'b1;
    assign upc_loop_intf_3.finish = finish;
    csv_file_dump upc_loop_csv_dumper_3;
    upc_loop_monitor #(2) upc_loop_monitor_3;
    upc_loop_intf#(2) upc_loop_intf_4(clock,reset);
    assign upc_loop_intf_4.cur_state = AESL_inst_dut.grp_dut_Pipeline_VITIS_LOOP_14_1_fu_5406.ap_CS_fsm;
    assign upc_loop_intf_4.iter_start_state = AESL_inst_dut.grp_dut_Pipeline_VITIS_LOOP_14_1_fu_5406.ap_ST_fsm_pp0_stage0;
    assign upc_loop_intf_4.iter_end_state = AESL_inst_dut.grp_dut_Pipeline_VITIS_LOOP_14_1_fu_5406.ap_ST_fsm_pp0_stage0;
    assign upc_loop_intf_4.quit_state = AESL_inst_dut.grp_dut_Pipeline_VITIS_LOOP_14_1_fu_5406.ap_ST_fsm_pp0_stage0;
    assign upc_loop_intf_4.iter_start_block = AESL_inst_dut.grp_dut_Pipeline_VITIS_LOOP_14_1_fu_5406.ap_block_pp0_stage0_subdone;
    assign upc_loop_intf_4.iter_end_block = AESL_inst_dut.grp_dut_Pipeline_VITIS_LOOP_14_1_fu_5406.ap_block_pp0_stage0_subdone;
    assign upc_loop_intf_4.quit_block = AESL_inst_dut.grp_dut_Pipeline_VITIS_LOOP_14_1_fu_5406.ap_block_pp0_stage0_subdone;
    assign upc_loop_intf_4.iter_start_enable = AESL_inst_dut.grp_dut_Pipeline_VITIS_LOOP_14_1_fu_5406.ap_enable_reg_pp0_iter0;
    assign upc_loop_intf_4.iter_end_enable = AESL_inst_dut.grp_dut_Pipeline_VITIS_LOOP_14_1_fu_5406.ap_enable_reg_pp0_iter1;
    assign upc_loop_intf_4.quit_enable = AESL_inst_dut.grp_dut_Pipeline_VITIS_LOOP_14_1_fu_5406.ap_enable_reg_pp0_iter1;
    assign upc_loop_intf_4.loop_start = AESL_inst_dut.grp_dut_Pipeline_VITIS_LOOP_14_1_fu_5406.ap_start;
    assign upc_loop_intf_4.loop_ready = AESL_inst_dut.grp_dut_Pipeline_VITIS_LOOP_14_1_fu_5406.ap_ready;
    assign upc_loop_intf_4.loop_done = AESL_inst_dut.grp_dut_Pipeline_VITIS_LOOP_14_1_fu_5406.ap_done_int;
    assign upc_loop_intf_4.loop_continue = 1'b1;
    assign upc_loop_intf_4.quit_at_end = 1'b1;
    assign upc_loop_intf_4.finish = finish;
    csv_file_dump upc_loop_csv_dumper_4;
    upc_loop_monitor #(2) upc_loop_monitor_4;
    upc_loop_intf#(1) upc_loop_intf_5(clock,reset);
    assign upc_loop_intf_5.cur_state = AESL_inst_dut.grp_divide_fu_5412.grp_divide_Pipeline_NORMALIZE_fu_2815.ap_CS_fsm;
    assign upc_loop_intf_5.iter_start_state = AESL_inst_dut.grp_divide_fu_5412.grp_divide_Pipeline_NORMALIZE_fu_2815.ap_ST_fsm_pp0_stage0;
    assign upc_loop_intf_5.iter_end_state = AESL_inst_dut.grp_divide_fu_5412.grp_divide_Pipeline_NORMALIZE_fu_2815.ap_ST_fsm_pp0_stage0;
    assign upc_loop_intf_5.quit_state = AESL_inst_dut.grp_divide_fu_5412.grp_divide_Pipeline_NORMALIZE_fu_2815.ap_ST_fsm_pp0_stage0;
    assign upc_loop_intf_5.iter_start_block = AESL_inst_dut.grp_divide_fu_5412.grp_divide_Pipeline_NORMALIZE_fu_2815.ap_block_pp0_stage0_subdone;
    assign upc_loop_intf_5.iter_end_block = AESL_inst_dut.grp_divide_fu_5412.grp_divide_Pipeline_NORMALIZE_fu_2815.ap_block_pp0_stage0_subdone;
    assign upc_loop_intf_5.quit_block = AESL_inst_dut.grp_divide_fu_5412.grp_divide_Pipeline_NORMALIZE_fu_2815.ap_block_pp0_stage0_subdone;
    assign upc_loop_intf_5.iter_start_enable = AESL_inst_dut.grp_divide_fu_5412.grp_divide_Pipeline_NORMALIZE_fu_2815.ap_enable_reg_pp0_iter1;
    assign upc_loop_intf_5.iter_end_enable = AESL_inst_dut.grp_divide_fu_5412.grp_divide_Pipeline_NORMALIZE_fu_2815.ap_enable_reg_pp0_iter1;
    assign upc_loop_intf_5.quit_enable = AESL_inst_dut.grp_divide_fu_5412.grp_divide_Pipeline_NORMALIZE_fu_2815.ap_enable_reg_pp0_iter1;
    assign upc_loop_intf_5.loop_start = AESL_inst_dut.grp_divide_fu_5412.grp_divide_Pipeline_NORMALIZE_fu_2815.ap_start;
    assign upc_loop_intf_5.loop_ready = AESL_inst_dut.grp_divide_fu_5412.grp_divide_Pipeline_NORMALIZE_fu_2815.ap_ready;
    assign upc_loop_intf_5.loop_done = AESL_inst_dut.grp_divide_fu_5412.grp_divide_Pipeline_NORMALIZE_fu_2815.ap_done_int;
    assign upc_loop_intf_5.loop_continue = 1'b1;
    assign upc_loop_intf_5.quit_at_end = 1'b1;
    assign upc_loop_intf_5.finish = finish;
    csv_file_dump upc_loop_csv_dumper_5;
    upc_loop_monitor #(1) upc_loop_monitor_5;
    upc_loop_intf#(2) upc_loop_intf_6(clock,reset);
    assign upc_loop_intf_6.cur_state = AESL_inst_dut.grp_divide_fu_5412.grp_divide_Pipeline_ADJUST_fu_2889.ap_CS_fsm;
    assign upc_loop_intf_6.iter_start_state = AESL_inst_dut.grp_divide_fu_5412.grp_divide_Pipeline_ADJUST_fu_2889.ap_ST_fsm_pp0_stage0;
    assign upc_loop_intf_6.iter_end_state = AESL_inst_dut.grp_divide_fu_5412.grp_divide_Pipeline_ADJUST_fu_2889.ap_ST_fsm_pp0_stage1;
    assign upc_loop_intf_6.quit_state = AESL_inst_dut.grp_divide_fu_5412.grp_divide_Pipeline_ADJUST_fu_2889.ap_ST_fsm_pp0_stage1;
    assign upc_loop_intf_6.iter_start_block = AESL_inst_dut.grp_divide_fu_5412.grp_divide_Pipeline_ADJUST_fu_2889.ap_block_pp0_stage0_subdone;
    assign upc_loop_intf_6.iter_end_block = AESL_inst_dut.grp_divide_fu_5412.grp_divide_Pipeline_ADJUST_fu_2889.ap_block_pp0_stage1_subdone;
    assign upc_loop_intf_6.quit_block = AESL_inst_dut.grp_divide_fu_5412.grp_divide_Pipeline_ADJUST_fu_2889.ap_block_pp0_stage1_subdone;
    assign upc_loop_intf_6.iter_start_enable = AESL_inst_dut.grp_divide_fu_5412.grp_divide_Pipeline_ADJUST_fu_2889.ap_enable_reg_pp0_iter0;
    assign upc_loop_intf_6.iter_end_enable = AESL_inst_dut.grp_divide_fu_5412.grp_divide_Pipeline_ADJUST_fu_2889.ap_enable_reg_pp0_iter1;
    assign upc_loop_intf_6.quit_enable = AESL_inst_dut.grp_divide_fu_5412.grp_divide_Pipeline_ADJUST_fu_2889.ap_enable_reg_pp0_iter0;
    assign upc_loop_intf_6.loop_start = AESL_inst_dut.grp_divide_fu_5412.grp_divide_Pipeline_ADJUST_fu_2889.ap_start;
    assign upc_loop_intf_6.loop_ready = AESL_inst_dut.grp_divide_fu_5412.grp_divide_Pipeline_ADJUST_fu_2889.ap_ready;
    assign upc_loop_intf_6.loop_done = AESL_inst_dut.grp_divide_fu_5412.grp_divide_Pipeline_ADJUST_fu_2889.ap_done_int;
    assign upc_loop_intf_6.loop_continue = 1'b1;
    assign upc_loop_intf_6.quit_at_end = 1'b0;
    assign upc_loop_intf_6.finish = finish;
    csv_file_dump upc_loop_csv_dumper_6;
    upc_loop_monitor #(2) upc_loop_monitor_6;
    upc_loop_intf#(8) upc_loop_intf_7(clock,reset);
    assign upc_loop_intf_7.cur_state = AESL_inst_dut.grp_operator_mul_fu_5426.grp_operator_Pipeline_OUTER_INNER_fu_371.ap_CS_fsm;
    assign upc_loop_intf_7.iter_start_state = AESL_inst_dut.grp_operator_mul_fu_5426.grp_operator_Pipeline_OUTER_INNER_fu_371.ap_ST_fsm_pp0_stage0;
    assign upc_loop_intf_7.iter_end_state = AESL_inst_dut.grp_operator_mul_fu_5426.grp_operator_Pipeline_OUTER_INNER_fu_371.ap_ST_fsm_pp0_stage4;
    assign upc_loop_intf_7.quit_state = AESL_inst_dut.grp_operator_mul_fu_5426.grp_operator_Pipeline_OUTER_INNER_fu_371.ap_ST_fsm_pp0_stage4;
    assign upc_loop_intf_7.iter_start_block = AESL_inst_dut.grp_operator_mul_fu_5426.grp_operator_Pipeline_OUTER_INNER_fu_371.ap_block_pp0_stage0_subdone;
    assign upc_loop_intf_7.iter_end_block = AESL_inst_dut.grp_operator_mul_fu_5426.grp_operator_Pipeline_OUTER_INNER_fu_371.ap_block_pp0_stage4_subdone;
    assign upc_loop_intf_7.quit_block = AESL_inst_dut.grp_operator_mul_fu_5426.grp_operator_Pipeline_OUTER_INNER_fu_371.ap_block_pp0_stage4_subdone;
    assign upc_loop_intf_7.iter_start_enable = AESL_inst_dut.grp_operator_mul_fu_5426.grp_operator_Pipeline_OUTER_INNER_fu_371.ap_enable_reg_pp0_iter0;
    assign upc_loop_intf_7.iter_end_enable = AESL_inst_dut.grp_operator_mul_fu_5426.grp_operator_Pipeline_OUTER_INNER_fu_371.ap_enable_reg_pp0_iter1;
    assign upc_loop_intf_7.quit_enable = AESL_inst_dut.grp_operator_mul_fu_5426.grp_operator_Pipeline_OUTER_INNER_fu_371.ap_enable_reg_pp0_iter1;
    assign upc_loop_intf_7.loop_start = AESL_inst_dut.grp_operator_mul_fu_5426.grp_operator_Pipeline_OUTER_INNER_fu_371.ap_start;
    assign upc_loop_intf_7.loop_ready = AESL_inst_dut.grp_operator_mul_fu_5426.grp_operator_Pipeline_OUTER_INNER_fu_371.ap_ready;
    assign upc_loop_intf_7.loop_done = AESL_inst_dut.grp_operator_mul_fu_5426.grp_operator_Pipeline_OUTER_INNER_fu_371.ap_done_int;
    assign upc_loop_intf_7.loop_continue = 1'b1;
    assign upc_loop_intf_7.quit_at_end = 1'b1;
    assign upc_loop_intf_7.finish = finish;
    csv_file_dump upc_loop_csv_dumper_7;
    upc_loop_monitor #(8) upc_loop_monitor_7;
    upc_loop_intf#(8) upc_loop_intf_8(clock,reset);
    assign upc_loop_intf_8.cur_state = AESL_inst_dut.grp_operator_1_fu_5440.grp_operator_1_Pipeline_OUTER_INNER_fu_369.ap_CS_fsm;
    assign upc_loop_intf_8.iter_start_state = AESL_inst_dut.grp_operator_1_fu_5440.grp_operator_1_Pipeline_OUTER_INNER_fu_369.ap_ST_fsm_pp0_stage0;
    assign upc_loop_intf_8.iter_end_state = AESL_inst_dut.grp_operator_1_fu_5440.grp_operator_1_Pipeline_OUTER_INNER_fu_369.ap_ST_fsm_pp0_stage4;
    assign upc_loop_intf_8.quit_state = AESL_inst_dut.grp_operator_1_fu_5440.grp_operator_1_Pipeline_OUTER_INNER_fu_369.ap_ST_fsm_pp0_stage4;
    assign upc_loop_intf_8.iter_start_block = AESL_inst_dut.grp_operator_1_fu_5440.grp_operator_1_Pipeline_OUTER_INNER_fu_369.ap_block_pp0_stage0_subdone;
    assign upc_loop_intf_8.iter_end_block = AESL_inst_dut.grp_operator_1_fu_5440.grp_operator_1_Pipeline_OUTER_INNER_fu_369.ap_block_pp0_stage4_subdone;
    assign upc_loop_intf_8.quit_block = AESL_inst_dut.grp_operator_1_fu_5440.grp_operator_1_Pipeline_OUTER_INNER_fu_369.ap_block_pp0_stage4_subdone;
    assign upc_loop_intf_8.iter_start_enable = AESL_inst_dut.grp_operator_1_fu_5440.grp_operator_1_Pipeline_OUTER_INNER_fu_369.ap_enable_reg_pp0_iter0;
    assign upc_loop_intf_8.iter_end_enable = AESL_inst_dut.grp_operator_1_fu_5440.grp_operator_1_Pipeline_OUTER_INNER_fu_369.ap_enable_reg_pp0_iter1;
    assign upc_loop_intf_8.quit_enable = AESL_inst_dut.grp_operator_1_fu_5440.grp_operator_1_Pipeline_OUTER_INNER_fu_369.ap_enable_reg_pp0_iter1;
    assign upc_loop_intf_8.loop_start = AESL_inst_dut.grp_operator_1_fu_5440.grp_operator_1_Pipeline_OUTER_INNER_fu_369.ap_start;
    assign upc_loop_intf_8.loop_ready = AESL_inst_dut.grp_operator_1_fu_5440.grp_operator_1_Pipeline_OUTER_INNER_fu_369.ap_ready;
    assign upc_loop_intf_8.loop_done = AESL_inst_dut.grp_operator_1_fu_5440.grp_operator_1_Pipeline_OUTER_INNER_fu_369.ap_done_int;
    assign upc_loop_intf_8.loop_continue = 1'b1;
    assign upc_loop_intf_8.quit_at_end = 1'b1;
    assign upc_loop_intf_8.finish = finish;
    csv_file_dump upc_loop_csv_dumper_8;
    upc_loop_monitor #(8) upc_loop_monitor_8;
    upc_loop_intf#(2) upc_loop_intf_9(clock,reset);
    assign upc_loop_intf_9.cur_state = AESL_inst_dut.grp_dut_Pipeline_WRITE_LOOP_fu_5446.ap_CS_fsm;
    assign upc_loop_intf_9.iter_start_state = AESL_inst_dut.grp_dut_Pipeline_WRITE_LOOP_fu_5446.ap_ST_fsm_pp0_stage0;
    assign upc_loop_intf_9.iter_end_state = AESL_inst_dut.grp_dut_Pipeline_WRITE_LOOP_fu_5446.ap_ST_fsm_pp0_stage1;
    assign upc_loop_intf_9.quit_state = AESL_inst_dut.grp_dut_Pipeline_WRITE_LOOP_fu_5446.ap_ST_fsm_pp0_stage1;
    assign upc_loop_intf_9.iter_start_block = AESL_inst_dut.grp_dut_Pipeline_WRITE_LOOP_fu_5446.ap_block_pp0_stage0_subdone;
    assign upc_loop_intf_9.iter_end_block = AESL_inst_dut.grp_dut_Pipeline_WRITE_LOOP_fu_5446.ap_block_pp0_stage1_subdone;
    assign upc_loop_intf_9.quit_block = AESL_inst_dut.grp_dut_Pipeline_WRITE_LOOP_fu_5446.ap_block_pp0_stage1_subdone;
    assign upc_loop_intf_9.iter_start_enable = AESL_inst_dut.grp_dut_Pipeline_WRITE_LOOP_fu_5446.ap_enable_reg_pp0_iter0;
    assign upc_loop_intf_9.iter_end_enable = AESL_inst_dut.grp_dut_Pipeline_WRITE_LOOP_fu_5446.ap_enable_reg_pp0_iter1;
    assign upc_loop_intf_9.quit_enable = AESL_inst_dut.grp_dut_Pipeline_WRITE_LOOP_fu_5446.ap_enable_reg_pp0_iter1;
    assign upc_loop_intf_9.loop_start = AESL_inst_dut.grp_dut_Pipeline_WRITE_LOOP_fu_5446.ap_start;
    assign upc_loop_intf_9.loop_ready = AESL_inst_dut.grp_dut_Pipeline_WRITE_LOOP_fu_5446.ap_ready;
    assign upc_loop_intf_9.loop_done = AESL_inst_dut.grp_dut_Pipeline_WRITE_LOOP_fu_5446.ap_done_int;
    assign upc_loop_intf_9.loop_continue = 1'b1;
    assign upc_loop_intf_9.quit_at_end = 1'b1;
    assign upc_loop_intf_9.finish = finish;
    csv_file_dump upc_loop_csv_dumper_9;
    upc_loop_monitor #(2) upc_loop_monitor_9;

    sample_manager sample_manager_inst;

initial begin
    sample_manager_inst = new;



    mstatus_csv_dumper_1 = new("./module_status1.csv");
    module_monitor_1 = new(module_intf_1,mstatus_csv_dumper_1);
    mstatus_csv_dumper_2 = new("./module_status2.csv");
    module_monitor_2 = new(module_intf_2,mstatus_csv_dumper_2);
    mstatus_csv_dumper_3 = new("./module_status3.csv");
    module_monitor_3 = new(module_intf_3,mstatus_csv_dumper_3);
    mstatus_csv_dumper_4 = new("./module_status4.csv");
    module_monitor_4 = new(module_intf_4,mstatus_csv_dumper_4);
    mstatus_csv_dumper_5 = new("./module_status5.csv");
    module_monitor_5 = new(module_intf_5,mstatus_csv_dumper_5);
    mstatus_csv_dumper_6 = new("./module_status6.csv");
    module_monitor_6 = new(module_intf_6,mstatus_csv_dumper_6);
    mstatus_csv_dumper_7 = new("./module_status7.csv");
    module_monitor_7 = new(module_intf_7,mstatus_csv_dumper_7);
    mstatus_csv_dumper_8 = new("./module_status8.csv");
    module_monitor_8 = new(module_intf_8,mstatus_csv_dumper_8);
    mstatus_csv_dumper_9 = new("./module_status9.csv");
    module_monitor_9 = new(module_intf_9,mstatus_csv_dumper_9);
    mstatus_csv_dumper_10 = new("./module_status10.csv");
    module_monitor_10 = new(module_intf_10,mstatus_csv_dumper_10);
    mstatus_csv_dumper_11 = new("./module_status11.csv");
    module_monitor_11 = new(module_intf_11,mstatus_csv_dumper_11);
    mstatus_csv_dumper_12 = new("./module_status12.csv");
    module_monitor_12 = new(module_intf_12,mstatus_csv_dumper_12);
    mstatus_csv_dumper_13 = new("./module_status13.csv");
    module_monitor_13 = new(module_intf_13,mstatus_csv_dumper_13);
    mstatus_csv_dumper_14 = new("./module_status14.csv");
    module_monitor_14 = new(module_intf_14,mstatus_csv_dumper_14);
    mstatus_csv_dumper_15 = new("./module_status15.csv");
    module_monitor_15 = new(module_intf_15,mstatus_csv_dumper_15);
    mstatus_csv_dumper_16 = new("./module_status16.csv");
    module_monitor_16 = new(module_intf_16,mstatus_csv_dumper_16);
    mstatus_csv_dumper_17 = new("./module_status17.csv");
    module_monitor_17 = new(module_intf_17,mstatus_csv_dumper_17);
    mstatus_csv_dumper_18 = new("./module_status18.csv");
    module_monitor_18 = new(module_intf_18,mstatus_csv_dumper_18);
    mstatus_csv_dumper_19 = new("./module_status19.csv");
    module_monitor_19 = new(module_intf_19,mstatus_csv_dumper_19);
    mstatus_csv_dumper_20 = new("./module_status20.csv");
    module_monitor_20 = new(module_intf_20,mstatus_csv_dumper_20);
    mstatus_csv_dumper_21 = new("./module_status21.csv");
    module_monitor_21 = new(module_intf_21,mstatus_csv_dumper_21);
    mstatus_csv_dumper_22 = new("./module_status22.csv");
    module_monitor_22 = new(module_intf_22,mstatus_csv_dumper_22);

    pp_loop_csv_dumper_1 = new("./pp_loop_status1.csv");
    pp_loop_monitor_1 = new(pp_loop_intf_1,pp_loop_csv_dumper_1);
    pp_loop_csv_dumper_2 = new("./pp_loop_status2.csv");
    pp_loop_monitor_2 = new(pp_loop_intf_2,pp_loop_csv_dumper_2);
    pp_loop_csv_dumper_3 = new("./pp_loop_status3.csv");
    pp_loop_monitor_3 = new(pp_loop_intf_3,pp_loop_csv_dumper_3);


    seq_loop_csv_dumper_1 = new("./seq_loop_status1.csv");
    seq_loop_monitor_1 = new(seq_loop_intf_1,seq_loop_csv_dumper_1);
    seq_loop_csv_dumper_2 = new("./seq_loop_status2.csv");
    seq_loop_monitor_2 = new(seq_loop_intf_2,seq_loop_csv_dumper_2);
    seq_loop_csv_dumper_3 = new("./seq_loop_status3.csv");
    seq_loop_monitor_3 = new(seq_loop_intf_3,seq_loop_csv_dumper_3);
    seq_loop_csv_dumper_4 = new("./seq_loop_status4.csv");
    seq_loop_monitor_4 = new(seq_loop_intf_4,seq_loop_csv_dumper_4);
    seq_loop_csv_dumper_5 = new("./seq_loop_status5.csv");
    seq_loop_monitor_5 = new(seq_loop_intf_5,seq_loop_csv_dumper_5);

    upc_loop_csv_dumper_1 = new("./upc_loop_status1.csv");
    upc_loop_monitor_1 = new(upc_loop_intf_1,upc_loop_csv_dumper_1);
    upc_loop_csv_dumper_2 = new("./upc_loop_status2.csv");
    upc_loop_monitor_2 = new(upc_loop_intf_2,upc_loop_csv_dumper_2);
    upc_loop_csv_dumper_3 = new("./upc_loop_status3.csv");
    upc_loop_monitor_3 = new(upc_loop_intf_3,upc_loop_csv_dumper_3);
    upc_loop_csv_dumper_4 = new("./upc_loop_status4.csv");
    upc_loop_monitor_4 = new(upc_loop_intf_4,upc_loop_csv_dumper_4);
    upc_loop_csv_dumper_5 = new("./upc_loop_status5.csv");
    upc_loop_monitor_5 = new(upc_loop_intf_5,upc_loop_csv_dumper_5);
    upc_loop_csv_dumper_6 = new("./upc_loop_status6.csv");
    upc_loop_monitor_6 = new(upc_loop_intf_6,upc_loop_csv_dumper_6);
    upc_loop_csv_dumper_7 = new("./upc_loop_status7.csv");
    upc_loop_monitor_7 = new(upc_loop_intf_7,upc_loop_csv_dumper_7);
    upc_loop_csv_dumper_8 = new("./upc_loop_status8.csv");
    upc_loop_monitor_8 = new(upc_loop_intf_8,upc_loop_csv_dumper_8);
    upc_loop_csv_dumper_9 = new("./upc_loop_status9.csv");
    upc_loop_monitor_9 = new(upc_loop_intf_9,upc_loop_csv_dumper_9);

    sample_manager_inst.add_one_monitor(module_monitor_1);
    sample_manager_inst.add_one_monitor(module_monitor_2);
    sample_manager_inst.add_one_monitor(module_monitor_3);
    sample_manager_inst.add_one_monitor(module_monitor_4);
    sample_manager_inst.add_one_monitor(module_monitor_5);
    sample_manager_inst.add_one_monitor(module_monitor_6);
    sample_manager_inst.add_one_monitor(module_monitor_7);
    sample_manager_inst.add_one_monitor(module_monitor_8);
    sample_manager_inst.add_one_monitor(module_monitor_9);
    sample_manager_inst.add_one_monitor(module_monitor_10);
    sample_manager_inst.add_one_monitor(module_monitor_11);
    sample_manager_inst.add_one_monitor(module_monitor_12);
    sample_manager_inst.add_one_monitor(module_monitor_13);
    sample_manager_inst.add_one_monitor(module_monitor_14);
    sample_manager_inst.add_one_monitor(module_monitor_15);
    sample_manager_inst.add_one_monitor(module_monitor_16);
    sample_manager_inst.add_one_monitor(module_monitor_17);
    sample_manager_inst.add_one_monitor(module_monitor_18);
    sample_manager_inst.add_one_monitor(module_monitor_19);
    sample_manager_inst.add_one_monitor(module_monitor_20);
    sample_manager_inst.add_one_monitor(module_monitor_21);
    sample_manager_inst.add_one_monitor(module_monitor_22);
    sample_manager_inst.add_one_monitor(pp_loop_monitor_1);
    sample_manager_inst.add_one_monitor(pp_loop_monitor_2);
    sample_manager_inst.add_one_monitor(pp_loop_monitor_3);
    sample_manager_inst.add_one_monitor(seq_loop_monitor_1);
    sample_manager_inst.add_one_monitor(seq_loop_monitor_2);
    sample_manager_inst.add_one_monitor(seq_loop_monitor_3);
    sample_manager_inst.add_one_monitor(seq_loop_monitor_4);
    sample_manager_inst.add_one_monitor(seq_loop_monitor_5);
    sample_manager_inst.add_one_monitor(upc_loop_monitor_1);
    sample_manager_inst.add_one_monitor(upc_loop_monitor_2);
    sample_manager_inst.add_one_monitor(upc_loop_monitor_3);
    sample_manager_inst.add_one_monitor(upc_loop_monitor_4);
    sample_manager_inst.add_one_monitor(upc_loop_monitor_5);
    sample_manager_inst.add_one_monitor(upc_loop_monitor_6);
    sample_manager_inst.add_one_monitor(upc_loop_monitor_7);
    sample_manager_inst.add_one_monitor(upc_loop_monitor_8);
    sample_manager_inst.add_one_monitor(upc_loop_monitor_9);
    
    fork
        sample_manager_inst.start_monitor();
        last_transaction_done;
    join
    disable fork;

    sample_manager_inst.start_dump();
end

    task last_transaction_done();
        wait(reset == 0);
        while(1) begin
            if (finish == 1'b1)
                break;
            else
                @(posedge clock);
        end
    endtask


endmodule
